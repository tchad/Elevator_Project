library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity INPUT_MUX is
  Port ( );
end INPUT_MUX;

architecture Behavioral of INPUT_MUX is

begin


end Behavioral;
